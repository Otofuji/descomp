library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity atividade1aula2 is
   generic (
          dataWidth: natural := 8;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture eric of atividade1aula2 is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
        -- Inicializa os endereços:
        tmp(0) := x"45";
        tmp(1) := x"52";
        tmp(2) := x"49";
        tmp(3) := x"43";
        tmp(4) := x"00";
        tmp(5) := x"10";
        tmp(6) := x"13";
        tmp(7) := x"12";
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;